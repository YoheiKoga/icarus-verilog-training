`timescale 1ns / 1ns
module stimulus();
    // input
    reg x;

endmodule // stimulus